interface axi_intf(input logic aclk, arst);


endinterface
