module axi_assertion();


endmodule
